module flatbuffers

pub fn decode<T>(b []byte) ?T {
	error('not implemented')
}
