module flatbuffers

pub fn encode<T>(object T) ?[]byte {
	error("not implemented")
}

struct VTable {
}

struct Table {
}

